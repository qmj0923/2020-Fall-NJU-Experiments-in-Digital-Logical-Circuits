module decoder_7seg(X, Y);
	input [3:0] X;
	output [6:0]Y;
	
	assign Y[0] = (X[3] & X[2] & X[1] & ~X[0]) | (X[3] & ~X[2] & X[1] & X[0]) | (~X[3] & X[2] & ~X[1] & ~X[0]) | (~X[3] & ~X[2] & X[1] & ~X[0]);
	
	assign Y[1] = (X[3] & ~X[2] & X[1] & ~X[0]) | (~X[2] & ~X[1] & X[0]) | (~X[3] & ~X[1] & ~X[0]) | (~X[3] & ~X[2] & X[0]);
	
	assign Y[2] = (X[3] & X[2] & ~X[1] & X[0]) | (~X[3] & ~X[2] & X[0]) | (~X[3] & ~X[2] & ~X[1]);
	
	assign Y[3] = (X[3] & X[2] & X[1] & ~X[0]) | (X[3] & ~X[2] & X[1] & X[0]) | (~X[2] & ~X[1] & ~X[0]) | (~X[3] & X[2] & ~X[1] & X[0]);
	
	assign Y[4] = (X[3] & ~X[0]) | (X[2] & X[1] & ~X[0]) | (X[3] & ~X[2] & X[1]);
	
	assign Y[5] = (X[3] & X[2] & ~X[0]) | (X[3] & X[2] & ~X[1]) | (X[3] & ~X[1] & ~X[0]) | (~X[3] & ~X[2] & X[1] & ~X[0]);
	
	assign Y[6] = (X[3] & X[2] & X[1]) | (X[3] & ~X[2] & ~X[1] & ~X[0]) | (~X[3] & ~X[2] & X[1] & X[0]);

endmodule 